-------------------------------------------------
-- Project : SPI Loopback      	              --
-- Author : Emiliano Sisinni                   --
-- Date : AY2022/2023                          --
-- Company : UniBS                             --
-- File : top_spiloopback.vhd                  --
-------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
--Assegnamento PIN FISICI
entity top_spiir is
	port(
		FPGA_CLK1_50: in std_logic;
		SW: in std_logic_vector(3 downto 0);
		KEY: in std_logic_vector(2 downto 0);
		LED: out std_logic_vector(1 downto 0);
		--PB: in std_logic_vector(1 downto 0);
		ARDUINO_IO: inout std_logic_vector(15 downto 0));
end top_spiir;

architecture top_arch of top_spiir is
begin

	spi0:entity work.basic_iir 
	generic map(
			DATA_W 	=> 16,			-- FIFO and SPI data width in bits
			Nbit 	=> 4 					-- log2(data width)
			)
	port map(
		OSC_FPGA => FPGA_CLK1_50,
		reset => '0',
		SYS_SPI_MOSI => ARDUINO_IO(11),--mosi
		SYS_SPI_MISO => ARDUINO_IO(12),
		SYS_SPI_SCK => ARDUINO_IO(13),
		LED => LED(1 downto 0)
		
		);
		
		ARDUINO_IO(7) <= ARDUINO_IO(11);--mosi
		ARDUINO_IO(6) <= ARDUINO_IO(12);--miso
		ARDUINO_IO(5) <= ARDUINO_IO(13);--sck
		

end top_arch;
